/*******************************************************************************
swankmania_HDL
Stephen Niedzielski - sniedzie@digipen.edu
*******************************************************************************/

`include "Global.h"

// Sony ACX705AKM controller.
// Created:   Friday, October 5, 2007 [Stephen Niedzielski]
// Modified:  Friday, October 5, 2007 [Stephen Niedzielski]
module ACX705AKM_Ctrl
(
  input         iClk100,
  input         iClk16,
  output        oVsync,
  output        oHsync,
  output        oSD,
  output        oMCK,  
  output [15:0] oAdr
);

  // Never shut down.
  assign oSD = 1'b1;

  localparam
  MCK_Hz        = 4_000_000,
  Hsync_Frame   = 200,
  Vsync_Hz      = 74, // ~74.171
  Dots_Frame    = 272,
  Pixels_Line   = 240,
  Lines_Frame   = 160,
  Pixels_Frame  = Pixels_Line * Lines_Frame;

  // Generate the 4 MHz MCK clock signal from a 16 MHz clock and two flip flops.
  reg
  _MCK8,
  _MCK;
  initial
  begin
    _MCK8 = 1'b0;
    _MCK = 1'b0;
  end
  assign oMCK = _MCK;

  // 16 MHz to 8 Mhz.
  always_ff @( posedge iClk16 )
  begin
    _MCK8 <= ~_MCK8;
  end

  // 8 Mhz to 4 MHz.
  always_ff @( posedge _MCK8 )
  begin
    _MCK <= ~_MCK;
  end
  
  reg
  _MCK100a,
  _MCK100b,
  _MCK100;
  initial
  begin
  _MCK100a = 1'bx;
  _MCK100b = 1'bx;
  _MCK100 = 1'bx;
  end
  
  wire MCK100;
  Debounce
  Debounce0
  (
    .iClk( iClk100 ),
    .iD( _MCK100 ),
    .oQ( MCK100 )
  );

  // HSYNC, VSYNC, and pixel management.
  reg [8:0] _DotCnt;
  reg [7:0] _HsyncCnt;
  initial
  begin
    _DotCnt = 9'h000;
    _HsyncCnt = 8'h00;
  end
  //assign oAdr = _DotCnt + Pixels_Line * _HsyncCnt;

  reg [8:0] _DotCnt100;
  reg [7:0] _HsyncCnt100;
  initial
  begin
    _DotCnt100 = 9'h000;
    _HsyncCnt100 = 8'h00;
  end
  assign oAdr = _DotCnt100 + Pixels_Line * _HsyncCnt100;

  // Dot count.
  always_ff @( posedge oMCK )
  begin
    if( _DotCnt == (Dots_Frame - 1'd1) )
      _DotCnt <= 9'h0;
    else
      _DotCnt <= _DotCnt + 1'd1;
  end
  
  reg _MCK100Dly;
  initial _MCK100Dly = 0;
  always_ff @( posedge iClk100 )
  begin
    _MCK100a <= _MCK;
    _MCK100b <= _MCK100a;
    _MCK100  <= _MCK100b;
    _MCK100Dly <= MCK100;
    
    if( MCK100 )
    begin
      if( _DotCnt100 == (Dots_Frame - 1'd1) )
        _DotCnt100 <= 9'h0;
      else
        _DotCnt100 <= _DotCnt100 + 1'd1;
    end
  end
  
  // Hsync count.
  always_ff @( posedge oMCK )
  begin
    if( _DotCnt == (Dots_Frame - 1'd1) )
    begin
      if( _HsyncCnt == (Hsync_Frame - 1'd1) )
        _HsyncCnt <= 8'h0;
      else
        _HsyncCnt <= _HsyncCnt + 1'd1;
    end
  end

  always_ff @( posedge iClk100 )
  begin
    if( _MCK100Dly && _DotCnt100 == (Dots_Frame - 1'd1) )
    begin
      if( _HsyncCnt100 == (Hsync_Frame - 1'd1) )
        _HsyncCnt100 <= 8'h0;
      else
        _HsyncCnt100 <= _HsyncCnt100 + 1'd1;
    end
  end
  
  // Hsync and Vsync.
  reg
  _Hsync,
  _Vsync;
  initial
  begin
    _Hsync = 1'b1;
    _Vsync = 1'b1;
  end
  always_ff @( posedge oMCK )
  begin
    // Note memory latency when outputting Vsync and Hsync.
    _Hsync <= _DotCnt >= 255 && _DotCnt <= 264 ? 1'b0 : 1'b1;
    _Vsync <= _HsyncCnt >= 180 && _HsyncCnt <= 182 ? 1'b0 : 1'b1;
  end
  assign
  oHsync = _Hsync,
  oVsync = _Vsync;

endmodule
